`timescale 1 ns / 1 ps

`include "ram.sv"
`include "decoder.sv"






