`timescale 1ns / 1ps
module alu_testbench;
    //Inputs
    reg[15:0] A,B;
    reg[3:0] ALU_Sel;
    //Outputs
    wire[15:0] ALU_Out;
    
endmodule